module nes6502(

);

endmodule